module prim_flop (
        clk_i,
        rst_ni,
        d_i,
        q_o
);
        parameter signed [31:0] Width = 1;
        parameter [Width - 1:0] ResetValue = 0;
        input clk_i;
        input rst_ni;
        input [Width - 1:0] d_i;
        output reg [Width - 1:0] q_o;
        always @(posedge clk_i or negedge rst_ni)
                if (!rst_ni)
                        q_o <= ResetValue;
                else
                        q_o <= d_i;
endmodule
